module sprite_rom (
	input [10:0]	addr,
	output [31:0]	data
);

	parameter ADDR_WIDTH = 11;
   parameter DATA_WIDTH =  8;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
		32'b00000000000000000000000000000000,
	};
	assign data = ROM[addr];
endmodule